library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity memoria_char is
port(
 addr : in std_logic_vector(10 downto 0);
 do : out std_logic_vector(7 downto 0)
 );
end memoria_char;

architecture syn of memoria_char is
type char_mem is array (0 to 1791) of std_logic_vector(7 downto 0);
constant char_ROM : char_mem := ( 
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+00 (nul)
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+01
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+02
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+03
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+04
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+05
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+06
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+07
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+08
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+09
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+0A
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+0B
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+0C
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+0D
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+0E
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+0F
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+10
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+11
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+12
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+13
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+14
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+15
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+16
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+17
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+18
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+19
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+1A
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+1B
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+1C
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+1D
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+1E
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+1F
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+20 (space)
     x"18", x"3C", x"3C", x"18", x"18", x"00", x"18", x"00",   -- U+21 (!)
     x"36", x"36", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+22 ()
     x"36", x"36", x"7F", x"36", x"7F", x"36", x"36", x"00",   -- U+23 (#)
     x"0C", x"3E", x"03", x"1E", x"30", x"1F", x"0C", x"00",   -- U+24 ($)
     x"00", x"63", x"33", x"18", x"0C", x"66", x"63", x"00",   -- U+25 (%)
     x"1C", x"36", x"1C", x"6E", x"3B", x"33", x"6E", x"00",   -- U+26 (&)
     x"06", x"06", x"03", x"00", x"00", x"00", x"00", x"00",   -- U+27 (')
     x"18", x"0C", x"06", x"06", x"06", x"0C", x"18", x"00",   -- U+28 (()
     x"06", x"0C", x"18", x"18", x"18", x"0C", x"06", x"00",   -- U+29 ())
     x"00", x"66", x"3C", x"FF", x"3C", x"66", x"00", x"00",   -- U+2A (*)
     x"00", x"0C", x"0C", x"3F", x"0C", x"0C", x"00", x"00",   -- U+2B (+)
     x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"06",   -- U+2C (,)
     x"00", x"00", x"00", x"3F", x"00", x"00", x"00", x"00",   -- U+2D (-)
     x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00",   -- U+2E (.)
     x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"00",   -- U+2F (/)
     x"3E", x"63", x"73", x"7B", x"6F", x"67", x"3E", x"00",   -- U+30 (0)
     x"0C", x"0E", x"0C", x"0C", x"0C", x"0C", x"3F", x"00",   -- U+31 (1)
     x"1E", x"33", x"30", x"1C", x"06", x"33", x"3F", x"00",   -- U+32 (2)
     x"1E", x"33", x"30", x"1C", x"30", x"33", x"1E", x"00",   -- U+33 (3)
     x"38", x"3C", x"36", x"33", x"7F", x"30", x"78", x"00",   -- U+34 (4)
     x"3F", x"03", x"1F", x"30", x"30", x"33", x"1E", x"00",   -- U+35 (5)
     x"1C", x"06", x"03", x"1F", x"33", x"33", x"1E", x"00",   -- U+36 (6)
     x"3F", x"33", x"30", x"18", x"0C", x"0C", x"0C", x"00",   -- U+37 (7)
     x"1E", x"33", x"33", x"1E", x"33", x"33", x"1E", x"00",   -- U+38 (8)
     x"1E", x"33", x"33", x"3E", x"30", x"18", x"0E", x"00",   -- U+39 (9)
     x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00",   -- U+3A (:)
     x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"06",   -- U+3B (;)
     x"18", x"0C", x"06", x"03", x"06", x"0C", x"18", x"00",   -- U+3C (<)
     x"00", x"00", x"3F", x"00", x"00", x"3F", x"00", x"00",   -- U+3D (=)
     x"06", x"0C", x"18", x"30", x"18", x"0C", x"06", x"00",   -- U+3E (>)
     x"1E", x"33", x"30", x"18", x"0C", x"00", x"0C", x"00",   -- U+3F (?)
     x"3E", x"63", x"7B", x"7B", x"7B", x"03", x"1E", x"00",   -- U+40 (@)
     x"0C", x"1E", x"33", x"33", x"3F", x"33", x"33", x"00",   -- U+41 (A)
     x"3F", x"66", x"66", x"3E", x"66", x"66", x"3F", x"00",   -- U+42 (B)
     x"3C", x"66", x"03", x"03", x"03", x"66", x"3C", x"00",   -- U+43 (C)
     x"1F", x"36", x"66", x"66", x"66", x"36", x"1F", x"00",   -- U+44 (D)
     x"7F", x"46", x"16", x"1E", x"16", x"46", x"7F", x"00",   -- U+45 (E)
     x"7F", x"46", x"16", x"1E", x"16", x"06", x"0F", x"00",   -- U+46 (F)
     x"3C", x"66", x"03", x"03", x"73", x"66", x"7C", x"00",   -- U+47 (G)
     x"33", x"33", x"33", x"3F", x"33", x"33", x"33", x"00",   -- U+48 (H)
     x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",   -- U+49 (I)
     x"78", x"30", x"30", x"30", x"33", x"33", x"1E", x"00",   -- U+4A (J)
     x"67", x"66", x"36", x"1E", x"36", x"66", x"67", x"00",   -- U+4B (K)
     x"0F", x"06", x"06", x"06", x"46", x"66", x"7F", x"00",   -- U+4C (L)
     x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",   -- U+4D (M)
     x"63", x"67", x"6F", x"7B", x"73", x"63", x"63", x"00",   -- U+4E (N)
     x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00",   -- U+4F (O)
     x"3F", x"66", x"66", x"3E", x"06", x"06", x"0F", x"00",   -- U+50 (P)
     x"1E", x"33", x"33", x"33", x"3B", x"1E", x"38", x"00",   -- U+51 (Q)
     x"3F", x"66", x"66", x"3E", x"36", x"66", x"67", x"00",   -- U+52 (R)
     x"1E", x"33", x"07", x"0E", x"38", x"33", x"1E", x"00",   -- U+53 (S)
     x"3F", x"2D", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",   -- U+54 (T)
     x"33", x"33", x"33", x"33", x"33", x"33", x"3F", x"00",   -- U+55 (U)
     x"33", x"33", x"33", x"33", x"33", x"1E", x"0C", x"00",   -- U+56 (V)
     x"63", x"63", x"63", x"6B", x"7F", x"77", x"63", x"00",   -- U+57 (W)
     x"63", x"63", x"36", x"1C", x"1C", x"36", x"63", x"00",   -- U+58 (X)
     x"33", x"33", x"33", x"1E", x"0C", x"0C", x"1E", x"00",   -- U+59 (Y)
     x"7F", x"63", x"31", x"18", x"4C", x"66", x"7F", x"00",   -- U+5A (Z)
     x"1E", x"06", x"06", x"06", x"06", x"06", x"1E", x"00",   -- U+5B ([)
     x"03", x"06", x"0C", x"18", x"30", x"60", x"40", x"00",   -- U+5C (\)
     x"1E", x"18", x"18", x"18", x"18", x"18", x"1E", x"00",   -- U+5D (])
     x"08", x"1C", x"36", x"63", x"00", x"00", x"00", x"00",   -- U+5E (^)
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",   -- U+5F (_)
     x"0C", x"0C", x"18", x"00", x"00", x"00", x"00", x"00",   -- U+60 (`)
     x"00", x"00", x"1E", x"30", x"3E", x"33", x"6E", x"00",   -- U+61 (a)
     x"07", x"06", x"06", x"3E", x"66", x"66", x"3B", x"00",   -- U+62 (b)
     x"00", x"00", x"1E", x"33", x"03", x"33", x"1E", x"00",   -- U+63 (c)
     x"38", x"30", x"30", x"3E", x"33", x"33", x"6E", x"00",   -- U+64 (d)
     x"00", x"00", x"1E", x"33", x"3F", x"03", x"1E", x"00",   -- U+65 (e)
     x"1C", x"36", x"06", x"0F", x"06", x"06", x"0F", x"00",   -- U+66 (f)
     x"00", x"00", x"6E", x"33", x"33", x"3E", x"30", x"1F",   -- U+67 (g)
     x"07", x"06", x"36", x"6E", x"66", x"66", x"67", x"00",   -- U+68 (h)
     x"0C", x"00", x"0E", x"0C", x"0C", x"0C", x"1E", x"00",   -- U+69 (i)
     x"30", x"00", x"30", x"30", x"30", x"33", x"33", x"1E",   -- U+6A (j)
     x"07", x"06", x"66", x"36", x"1E", x"36", x"67", x"00",   -- U+6B (k)
     x"0E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00",   -- U+6C (l)
     x"00", x"00", x"33", x"7F", x"7F", x"6B", x"63", x"00",   -- U+6D (m)
     x"00", x"00", x"1F", x"33", x"33", x"33", x"33", x"00",   -- U+6E (n)
     x"00", x"00", x"1E", x"33", x"33", x"33", x"1E", x"00",   -- U+6F (o)
     x"00", x"00", x"3B", x"66", x"66", x"3E", x"06", x"0F",   -- U+70 (p)
     x"00", x"00", x"6E", x"33", x"33", x"3E", x"30", x"78",   -- U+71 (q)
     x"00", x"00", x"3B", x"6E", x"66", x"06", x"0F", x"00",   -- U+72 (r)
     x"00", x"00", x"3E", x"03", x"1E", x"30", x"1F", x"00",   -- U+73 (s)
     x"08", x"0C", x"3E", x"0C", x"0C", x"2C", x"18", x"00",   -- U+74 (t)
     x"00", x"00", x"33", x"33", x"33", x"33", x"6E", x"00",   -- U+75 (u)
     x"00", x"00", x"33", x"33", x"33", x"1E", x"0C", x"00",   -- U+76 (v)
     x"00", x"00", x"63", x"6B", x"7F", x"7F", x"36", x"00",   -- U+77 (w)
     x"00", x"00", x"63", x"36", x"1C", x"36", x"63", x"00",   -- U+78 (x)
     x"00", x"00", x"33", x"33", x"33", x"3E", x"30", x"1F",   -- U+79 (y)
     x"00", x"00", x"3F", x"19", x"0C", x"26", x"3F", x"00",   -- U+7A (z)
     x"38", x"0C", x"0C", x"07", x"0C", x"0C", x"38", x"00",   -- U+7B ({)
     x"18", x"18", x"18", x"00", x"18", x"18", x"18", x"00",   -- U+7C (|)
     x"07", x"0C", x"0C", x"38", x"0C", x"0C", x"07", x"00",   -- U+7D (})
     x"6E", x"3B", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+7E (~)
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+7F
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+A0 (no break space)
     x"18", x"18", x"00", x"18", x"18", x"18", x"18", x"00",   -- U+A1 (inverted !)
     x"18", x"18", x"7E", x"03", x"03", x"7E", x"18", x"18",   -- U+A2 (dollarcents)
     x"1C", x"36", x"26", x"0F", x"06", x"67", x"3F", x"00",   -- U+A3 (pound sterling)
     x"00", x"00", x"63", x"3E", x"36", x"3E", x"63", x"00",   -- U+A4 (currency mark)
     x"33", x"33", x"1E", x"3F", x"0C", x"3F", x"0C", x"0C",   -- U+A5 (yen)
     x"18", x"18", x"18", x"00", x"18", x"18", x"18", x"00",   -- U+A6 (broken pipe)
     x"7C", x"C6", x"1C", x"36", x"36", x"1C", x"33", x"1E",   -- U+A7 (paragraph)
     x"33", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+A8 (diaeresis)
     x"3C", x"42", x"99", x"85", x"85", x"99", x"42", x"3C",   -- U+A9 (copyright symbol)
     x"3C", x"36", x"36", x"7C", x"00", x"00", x"00", x"00",   -- U+AA (superscript a)
     x"00", x"CC", x"66", x"33", x"66", x"CC", x"00", x"00",   -- U+AB (<<)
     x"00", x"00", x"00", x"3F", x"30", x"30", x"00", x"00",   -- U+AC (gun pointing left)
     x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+AD (soft hyphen)
     x"3C", x"42", x"9D", x"A5", x"9D", x"A5", x"42", x"3C",   -- U+AE (registered symbol)
     x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+AF (macron)
     x"1C", x"36", x"36", x"1C", x"00", x"00", x"00", x"00",   -- U+B0 (degree)
     x"18", x"18", x"7E", x"18", x"18", x"00", x"7E", x"00",   -- U+B1 (plusminus)
     x"1C", x"30", x"18", x"0C", x"3C", x"00", x"00", x"00",   -- U+B2 (superscript 2)
     x"1C", x"30", x"18", x"30", x"1C", x"00", x"00", x"00",   -- U+B2 (superscript 3)
     x"18", x"0C", x"00", x"00", x"00", x"00", x"00", x"00",   -- U+B2 (aigu)
     x"00", x"00", x"66", x"66", x"66", x"3E", x"06", x"03",   -- U+B5 (mu)
     x"FE", x"DB", x"DB", x"DE", x"D8", x"D8", x"D8", x"00",   -- U+B6 (pilcrow)
     x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00",   -- U+B7 (central dot)
     x"00", x"00", x"00", x"00", x"00", x"18", x"30", x"1E",   -- U+B8 (cedille)
     x"08", x"0C", x"08", x"1C", x"00", x"00", x"00", x"00",   -- U+B9 (superscript 1)
     x"1C", x"36", x"36", x"1C", x"00", x"00", x"00", x"00",   -- U+BA (superscript 0)
     x"00", x"33", x"66", x"CC", x"66", x"33", x"00", x"00",   -- U+BB (>>)
     x"C3", x"63", x"33", x"BD", x"EC", x"F6", x"F3", x"03",   -- U+BC (1/4)
     x"C3", x"63", x"33", x"7B", x"CC", x"66", x"33", x"F0",   -- U+BD (1/2)
     x"03", x"C4", x"63", x"B4", x"DB", x"AC", x"E6", x"80",   -- U+BE (3/4)
     x"0C", x"00", x"0C", x"06", x"03", x"33", x"1E", x"00",   -- U+BF (inverted ?)
     x"07", x"00", x"1C", x"36", x"63", x"7F", x"63", x"00",   -- U+C0 (A grave)
     x"70", x"00", x"1C", x"36", x"63", x"7F", x"63", x"00",   -- U+C1 (A aigu)
     x"1C", x"36", x"00", x"3E", x"63", x"7F", x"63", x"00",   -- U+C2 (A circumflex)
     x"6E", x"3B", x"00", x"3E", x"63", x"7F", x"63", x"00",   -- U+C3 (A ~)
     x"63", x"1C", x"36", x"63", x"7F", x"63", x"63", x"00",   -- U+C4 (A umlaut)
     x"0C", x"0C", x"00", x"1E", x"33", x"3F", x"33", x"00",   -- U+C5 (A ring)
     x"7C", x"36", x"33", x"7F", x"33", x"33", x"73", x"00",   -- U+C6 (AE)
     x"1E", x"33", x"03", x"33", x"1E", x"18", x"30", x"1E",   -- U+C7 (C cedille)
     x"07", x"00", x"3F", x"06", x"1E", x"06", x"3F", x"00",   -- U+C8 (E grave)
     x"38", x"00", x"3F", x"06", x"1E", x"06", x"3F", x"00",   -- U+C9 (E aigu)
     x"0C", x"12", x"3F", x"06", x"1E", x"06", x"3F", x"00",   -- U+CA (E circumflex)
     x"36", x"00", x"3F", x"06", x"1E", x"06", x"3F", x"00",   -- U+CB (E umlaut)
     x"07", x"00", x"1E", x"0C", x"0C", x"0C", x"1E", x"00",   -- U+CC (I grave)
     x"38", x"00", x"1E", x"0C", x"0C", x"0C", x"1E", x"00",   -- U+CD (I aigu)
     x"0C", x"12", x"00", x"1E", x"0C", x"0C", x"1E", x"00",   -- U+CE (I circumflex)
     x"33", x"00", x"1E", x"0C", x"0C", x"0C", x"1E", x"00",   -- U+CF (I umlaut)
     x"3F", x"66", x"6F", x"6F", x"66", x"66", x"3F", x"00",   -- U+D0 (Eth)
     x"3F", x"00", x"33", x"37", x"3F", x"3B", x"33", x"00",   -- U+D1 (N ~)
     x"0E", x"00", x"18", x"3C", x"66", x"3C", x"18", x"00",   -- U+D2 (O grave)
     x"70", x"00", x"18", x"3C", x"66", x"3C", x"18", x"00",   -- U+D3 (O aigu)
     x"3C", x"66", x"18", x"3C", x"66", x"3C", x"18", x"00",   -- U+D4 (O circumflex)
     x"6E", x"3B", x"00", x"3E", x"63", x"63", x"3E", x"00",   -- U+D5 (O ~)
     x"C3", x"18", x"3C", x"66", x"66", x"3C", x"18", x"00",   -- U+D6 (O umlaut)
     x"00", x"36", x"1C", x"08", x"1C", x"36", x"00", x"00",   -- U+D7 (multiplicative x)
     x"5C", x"36", x"73", x"7B", x"6F", x"36", x"1D", x"00",   -- U+D8 (O stroke)
     x"0E", x"00", x"66", x"66", x"66", x"66", x"3C", x"00",   -- U+D9 (U grave)
     x"70", x"00", x"66", x"66", x"66", x"66", x"3C", x"00",   -- U+DA (U aigu)
     x"3C", x"66", x"00", x"66", x"66", x"66", x"3C", x"00",   -- U+DB (U circumflex)
     x"33", x"00", x"33", x"33", x"33", x"33", x"1E", x"00",   -- U+DC (U umlaut)
     x"70", x"00", x"66", x"66", x"3C", x"18", x"18", x"00",   -- U+DD (Y aigu)
     x"0F", x"06", x"3E", x"66", x"66", x"3E", x"06", x"0F",   -- U+DE (Thorn)
     x"00", x"1E", x"33", x"1F", x"33", x"1F", x"03", x"03",   -- U+DF (beta)
     x"07", x"00", x"1E", x"30", x"3E", x"33", x"7E", x"00",   -- U+E0 (a grave)
     x"38", x"00", x"1E", x"30", x"3E", x"33", x"7E", x"00",   -- U+E1 (a aigu)
     x"7E", x"C3", x"3C", x"60", x"7C", x"66", x"FC", x"00",   -- U+E2 (a circumflex)
     x"6E", x"3B", x"1E", x"30", x"3E", x"33", x"7E", x"00",   -- U+E3 (a ~)
     x"33", x"00", x"1E", x"30", x"3E", x"33", x"7E", x"00",   -- U+E4 (a umlaut)
     x"0C", x"0C", x"1E", x"30", x"3E", x"33", x"7E", x"00",   -- U+E5 (a ring)
     x"00", x"00", x"FE", x"30", x"FE", x"33", x"FE", x"00",   -- U+E6 (ae)
     x"00", x"00", x"1E", x"03", x"03", x"1E", x"30", x"1C",   -- U+E7 (c cedille)
     x"07", x"00", x"1E", x"33", x"3F", x"03", x"1E", x"00",   -- U+E8 (e grave)
     x"38", x"00", x"1E", x"33", x"3F", x"03", x"1E", x"00",   -- U+E9 (e aigu)
     x"7E", x"C3", x"3C", x"66", x"7E", x"06", x"3C", x"00",   -- U+EA (e circumflex)
     x"33", x"00", x"1E", x"33", x"3F", x"03", x"1E", x"00",   -- U+EB (e umlaut)
     x"07", x"00", x"0E", x"0C", x"0C", x"0C", x"1E", x"00",   -- U+EC (i grave)
     x"1C", x"00", x"0E", x"0C", x"0C", x"0C", x"1E", x"00",   -- U+ED (i augu)
     x"3E", x"63", x"1C", x"18", x"18", x"18", x"3C", x"00",   -- U+EE (i circumflex)
     x"33", x"00", x"0E", x"0C", x"0C", x"0C", x"1E", x"00",   -- U+EF (i umlaut)
     x"1B", x"0E", x"1B", x"30", x"3E", x"33", x"1E", x"00",   -- U+F0 (eth)
     x"00", x"1F", x"00", x"1F", x"33", x"33", x"33", x"00",   -- U+F1 (n ~)
     x"00", x"07", x"00", x"1E", x"33", x"33", x"1E", x"00",   -- U+F2 (o grave)
     x"00", x"38", x"00", x"1E", x"33", x"33", x"1E", x"00",   -- U+F3 (o aigu)
     x"1E", x"33", x"00", x"1E", x"33", x"33", x"1E", x"00",   -- U+F4 (o circumflex)
     x"6E", x"3B", x"00", x"1E", x"33", x"33", x"1E", x"00",   -- U+F5 (o ~)
     x"00", x"33", x"00", x"1E", x"33", x"33", x"1E", x"00",   -- U+F6 (o umlaut)
     x"18", x"18", x"00", x"7E", x"00", x"18", x"18", x"00",   -- U+F7 (division)
     x"00", x"60", x"3C", x"76", x"7E", x"6E", x"3C", x"06",   -- U+F8 (o stroke)
     x"00", x"07", x"00", x"33", x"33", x"33", x"7E", x"00",   -- U+F9 (u grave)
     x"00", x"38", x"00", x"33", x"33", x"33", x"7E", x"00",   -- U+FA (u aigu)
     x"1E", x"33", x"00", x"33", x"33", x"33", x"7E", x"00",   -- U+FB (u circumflex)
     x"00", x"33", x"00", x"33", x"33", x"33", x"7E", x"00",   -- U+FC (u umlaut)
     x"00", x"38", x"00", x"33", x"33", x"3E", x"30", x"1F",   -- U+FD (y aigu)
     x"00", x"00", x"06", x"3E", x"66", x"3E", x"06", x"00",   -- U+FE (thorn)
     x"00", x"33", x"00", x"33", x"33", x"3E", x"30", x"1F");   -- U+FF (y umlaut)

begin

    do <= char_ROM(to_integer(unsigned(addr)));

end syn;